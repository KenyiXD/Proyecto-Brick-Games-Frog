LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY registro_universal_carros6 IS
	PORT(clock,reset,en,en2,R,L,enR,enL: IN STD_LOGIC;
		 Ent,Ent2: IN STD_LOGIC_VECTOR(7 downto 0);
		 Q : buffer STD_LOGIC_VECTOR (7 downto 0));
END registro_universal_carros6;

ARCHITECTURE solution OF registro_universal_carros6 IS

BEGIN
	PROCESS(clock,reset)
	BEGIN
		if reset='0' then Q<="10101010";
		elsif (clock'event and clock='1') then
			if(en='1') then 
				Q<=Ent;
			elsif(enR='1') then
				desplazamiento: for i in 6 downto 0 loop
				Q(i) <= Q(i+1);
				end loop;
				Q(7) <= R;
			elsif(enL='1') then
				desplazamiento1: for i in 1 to 7 loop  
                Q(i)<= Q(i-1);  
				end loop;  
				Q(0)<= L;
			elsif(en2='1') then
				Q<=Ent2;
			end if;
		end if;
	end process;
END solution;
